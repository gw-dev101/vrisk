module main

fn main() {
	println('Hello from vrisk!')
	println('This is a V project.')
}
