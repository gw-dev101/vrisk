module utils

// greet returns a greeting message for the given name
pub fn greet(name string) string {
	return 'Hello, ${name}! Welcome to vrisk.'
}

// add returns the sum of two integers
pub fn add(a int, b int) int {
	return a + b
}
